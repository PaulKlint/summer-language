# flex -- flexible arrays #

class flex ()
begin fetch update, retrieve, append, delete, size, next, 
            index, top;
      store size : change_size;

      var mem, size;

      proc extend()
      ( var i, m1 := array(mem.size + 10, undefined);
        for i in mem.index do m1[i] := mem[i] od;
        mem := m1
      );

      proc retrieve(i)
      if 0 <= i < size then return(mem[i]) else stop(-1) fi;

      proc update(i, v)
      if 0 <= i < size then return(mem[i] := v) else stop(-1) fi;

      proc append(v)
      ( if size >= mem.size then extend fi;
        mem[size] := v;
        size := size + 1;
        return(v)
      );

      proc delete(n)
      ( if size - n <= 0 then freturn else size := size - n fi );

      proc change_size(n)
      if n < 0 then freturn
      else
         if n >= mem.size then extend fi;
         return(size := n)
      fi;

      proc next(state)
      ( if state = undefined then state := 0 fi;
        if state < size then
           return([mem[state], state + 1])
        else
           freturn
        fi
      );

      proc index() return(interval(0, size - 1, 1));

      proc top()
      if size = 0 then freturn else return(mem[size-1]) fi;

init: mem := array(10, undefined);
      size := 0;
end flex;

var nstates := 0;
class item(name, body, dot, start, deriv)
begin fetch name, body, dot, start, deriv, focus, final,
            print, isterm, isnonterm, printderiv;
      
      proc focus()
        if dot < body.size then return(body[dot]) else freturn fi;

      proc final()
        return(dot = body.size);

      proc isterm()
        return((dot<body.size) & (body[dot] < 'A' | body[dot] > 'Z'));

      proc isnonterm()
        return((dot<body.size) & ('A' <= body[dot] <= 'Z'));

      proc print()
      ( var i;
        put('[', name, '->');
        for i in body.index
        do if i = dot then put('.') fi;
           put(body[i])
        od;
        if dot = body.size then put('.') fi;
        put(' , ', start, ']\n');
      );

      proc printderiv(indent)
      ( var d, pad2 := ' '.repl(indent+2);
	put(name, '->');
        if deriv.size = 1 & type(deriv[0]) = 'item' then
           deriv[0].printderiv(indent+2)
        else
           for d in deriv
           do case type(d) of
              'string':	put(d, ' '),
              'item':	put(d.name, ' ')
	      esac
	   od;
           put('\n');
           for d in deriv
           do if type(d) = 'item' then
                 put(pad2); d.printderiv(indent+2)
              fi
           od;
        fi
      );
init: nstates := nstates + 1;

end item;

class item_list()
begin fetch additem, next, print;
      var repr := flex;

      proc additem(name, body, dot, start, deriv, deriv_incr, look_ahead)
      ( var it, c;
	if dot < body.size & c := body[dot] &
	   (c < 'A' | c > 'Z') & c ~= look_ahead
	then
	   freturn
	fi;
        for it in repr
        do if it.name = name & it.body = body &
              it.dot = dot & it.start = start
           then
              freturn
           fi
        od;
	if deriv_incr ~= undefined
        then
           if deriv = undefined then
              deriv := flex
           elif type(deriv) = 'flex' then
              deriv := copy(deriv)
           elif type(deriv) = 'string' then
              deriv := flex.append(deriv)
           else
              put('deriv has illegal type'); stop(-1)
           fi;
           deriv.append(deriv_incr);
        fi;
        repr.append(item(name, body, dot, start, deriv));
        return
      );

      proc next(state) return(repr.next(state));

      proc print()
      ( var it;
        for it in repr do it.print od
      );

end item_list;

proc parse(P, start, inp)
( var A, B, I, j, p, change, n := inp.size, look_ahead := inp[0];

  I := array(n+1, undefined);
  for j in I.index do I[j] := item_list od;
  for p in P[start]
  do I[0].additem(start, p, 0, 0, undefined, undefined, look_ahead) | 'succeed' od;
  change := 1;
  while change ~= 0
  do change := 0;
     for B in I[0]
     do if B.final then
           for A in I[0]
           do if A.isnonterm & A.focus = B.name &
		 I[0].additem(A.name, A.body, A.dot+1, 0,
			      undefined, undefined, look_ahead) | 'succeed'
	      then
		 change := 1
              fi
           od
        fi
     od;
     for B in I[0]
     do if B.isnonterm then
           for p in P[B.focus]
           do if I[0].additem(B.focus, p, 0, 0, undefined, undefined, look_ahead) then
                 change := 1;
              fi
           od
        fi
     od;
  od;
  for j in interval(1, n, 1)
  do look_ahead := if j = n then undefined else inp[j] fi;
     for B in I[j-1]
     do					# scanner #
        if B.isterm & B.focus = inp[j-1] &
           I[j].additem(B.name, B.body, B.dot+1, B.start,
			B.deriv, inp[j-1], look_ahead)
	then # noop #
        fi;
     od;
     change := 1;
     while change ~= 0
     do change := 0;
        for A in I[j]
        do if A.final then		# completer #
              for B in I[A.start]
              do if B.isnonterm & B.focus = A.name &
                    I[j].additem(B.name, B.body, B.dot+1, B.start,
				 B.deriv, A, look_ahead)
                 then
                    change := 1;
                 fi;
              od;
           fi;
           if A.isnonterm then		# predictor #
              for p in P[A.focus]
              do if I[j].additem(A.focus, p, 0, j,
				 undefined, undefined, look_ahead) then
                    change := 1;
		 fi
              od
           fi
        od
     od;
   od;
   return(I);
);

proc do_parse(g, gname, startsymbol, phrase)
( var I, j, it ;
  nstates := 0;
  put('Parse "', phrase, '" with grammer "', gname, '"\n');
  I := parse(g, startsymbol, phrase);
#
  for j in I.index
  do put('I[', j, ']:\n');
     for it in I[j] do put('\t'); it.print od;
  od;
#
  put(nstates, ' states generated\n');
  for it in I[I.size-1]
  do if it.name = startsymbol & it.final & it.start = 0
     then put('Parse derived from: '); it.print;
          put('\n\n'); it.printderiv(0);
     fi;
  od;
);

var gram_ae :=
['E':	['T+E', 'T'],
 'T':	['F*T', 'F'],
 'F':	['(E)', 'a']
];
var sent_ae := ['(a+a)*a'];

var gram_ubda :=
['A':	['x', 'AA']];
var sent_ubda := ['xxxx'];

var gram_pal :=
['A':	['x', 'xAx']];
var sent_pal := ['xxxxx'];

var gram_gre :=
['X':	['a', 'Xb', 'Ya'],
 'Y':	['e', 'YdY']];
var sent_gre := ['ededea', 'ededeabbbb', 'ededededeabb'];

var gram_prop :=
['F':	['C', 'S', 'P', 'U'],
 'C':	['U>U'],
 'U':	['(F)', '~U', 'L'],
 'L':	['L`', 'p', 'q', 'r'],
 'S':	['U|S', 'U|U'],
 'P':	['U&P', 'U&U']];
var sent_prop :=
	[ 'p', '(p&q)', '(p`&q)|r|p|q`',
	  'p>((q>~(r`|(p&q)))>(q`|r))',
	  '~(~p`&(q|r)&p`)',
	  '((p&q)|(q&r)|(r&p`))>~((p`|q`)&(r`|p))'
	];

program early()
( var s;
  for s in sent_ae do do_parse(gram_ae, 'gram_ae', 'E', s) od;
  for s in sent_ubda do do_parse(gram_ubda, 'gram_ubda', 'A', s) od;
  for s in sent_pal do do_parse(gram_pal, 'gram_pal', 'A', s) od;
  for s in sent_gre do do_parse(gram_gre, 'gram_gre', 'X', s) od;
  for s in sent_prop do do_parse(gram_prop, 'gram_prop', 'F', s) od;
)
